
`define 	R_Type	7'b0110011
`define		Lw	7'b0000011
`define 	I_Type	7'b0010011
`define 	Jalr	7'b1100111
`define		J_Type	7'b1101111
`define		S_Type	7'b0100011
`define		U_Type	7'b0110111
`define 	B_Type	7'b1100011
`define 	Sub	10'b0100_0000_00
`define		Add	10'b0000_0000_00
`define 	Or	10'b0000_0001_10
`define		And	10'b0000_0001_11
`define		Sltu 10'b0000_0000_11
`define		Slt	10'b0000_0000_10
`define 	addi	3'b000
`define		lw	3'b010
`define 	ori	3'b110
`define		xori	3'b100
`define  	sltiu 3'b011
`define		slti	3'b010
`define		beq	3'b000
`define		jalr	3'b000
`define		blt	3'b100
`define 	bne	3'b001

`define 	bge	3'b101

module Controller(
	input[2:0] func3,
	input[6:0] func7,op,
	output reg MemWrite,ALUSrc,RegWrite,Jump,Branch,Jalr,
	output reg [1:0] ResultSrc,
	output reg [2:0] ALUControl,ImmSrc
	);


	wire[9:0] func;

	assign func={func7,func3};

	always@(func3,func7,op) begin

		{MemWrite,ALUSrc ,RegWrite,  Jump,Branch ,Jalr,ResultSrc,ALUControl ,ImmSrc}=14'b0000_0000_0100_00;
		case(op)

			`R_Type:begin

				RegWrite=1'b1;

				case(func)

					`Add: ALUControl=3'b010;
					`Sub:ALUControl=3'b110;
					`And:ALUControl =3'b000;
					`Or :ALUControl=3'b001;
					`Slt:ALUControl=3'b100;
					`Sltu:ALUControl= 3'b111;
				endcase

				end

			`Lw: {RegWrite ,ResultSrc, ALUSrc} = 4'b1011;

			`I_Type:begin

				{ ALUSrc, RegWrite } = 2'b11;
				case(func3)					
					`addi:ALUControl=3'b010;

					`xori:ALUControl=3'b011;
					`ori :ALUControl=3'b001;

					`slti:ALUControl=3'b100;

					`sltiu: begin ALUControl=3'b111; ImmSrc = 3'b101; end
				endcase
				end
			`Jalr:	{Jalr,ALUSrc, ResultSrc,RegWrite}=5'b11101;
			`S_Type:	{ImmSrc ,ALUSrc ,MemWrite}=5'b00111;

			`J_Type:	{ResultSrc, ImmSrc ,RegWrite, Jump}=7'b1001111;
			`B_Type:begin 

				{Branch,ImmSrc}=4'b1010;

				case(func3)

					`beq:	ALUControl=3'b110;
					`bne:	ALUControl=3'b110;

					`blt:	ALUControl=3'b111; 

					`bge:	ALUControl=3'b111;
				endcase
				end
				
			`U_Type:	{ResultSrc,ImmSrc,RegWrite}=6'b111001;
		endcase
	end
endmodule